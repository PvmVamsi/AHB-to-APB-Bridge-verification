package pkg;
	import uvm_pkg::*;
	
	`include "uvm_macros.svh"
	`include "mst_cfg.sv"
	`include "slv_cfg.sv"
	`include "env_cfg.sv"
	
	
	`include "mst_xtn.sv"
	`include "mst_seq.sv"
	`include "mst_seqr.sv"
	`include "mst_drv.sv"
	`include "mst_mon.sv"
	`include "mst_agt.sv"
	`include "mst_agt_top.sv"
	
	`include "slv_xtn.sv"
	`include "slv_seq.sv"
	`include "slv_seqr.sv"
	`include "slv_drv.sv"
	`include "slv_mon.sv"
	`include "slv_agt.sv"
	`include "slv_agt_top.sv"

	`include "vseqr.sv"
	`include "vseq.sv"
	`include "sb.sv"
	`include "env.sv"
	`include "test.sv"
endpackage
